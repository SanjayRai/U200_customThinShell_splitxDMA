// Year-Month-Date-Rev (YYMMDDVV)
`define SHELL_VERSION_NUMBER 32'h20083001
