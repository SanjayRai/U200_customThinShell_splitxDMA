// Sanjay Rai (sanjay.d.rai@gmail.com)
//
`timescale 1 ps / 1 ps

`include "shell_parameters.vh"

module shell_top (
  input [3:0]BMC_GPIO,
  input BMC_UART_rxd,
  output BMC_UART_txd,
  input C1_SYS_CLK,
  input [7:0]C0_DDR_SREF_CTRL_IN,
  output [7:0]C0_DDR_SREF_CTRL_OUT,
  input [7:0]C2_DDR_SREF_CTRL_IN,
  output [7:0]C2_DDR_SREF_CTRL_OUT,
  input [7:0]C3_DDR_SREF_CTRL_IN,
  output [7:0]C3_DDR_SREF_CTRL_OUT,
  hlx_AXI_LITE_intfc.master M_AXI_LITE_TO_HLS_PR_NORTH, 
  hlx_AXI_MM_intfc.slave S_AXI_MM_MIG, 
  hlx_AXI_MM_intfc.slave S_AXI_MM_PCIM, 
  output axi_reset_n_out,
  output c1_ddr4_act_n,
  output [16:0]c1_ddr4_adr,
  output [1:0]c1_ddr4_ba,
  output [1:0]c1_ddr4_bg,
  output [0:0]c1_ddr4_ck_c,
  output [0:0]c1_ddr4_ck_t,
  output [0:0]c1_ddr4_cke,
  output [0:0]c1_ddr4_cs_n,
  inout [71:0]c1_ddr4_dq,
  inout [17:0]c1_ddr4_dqs_c,
  inout [17:0]c1_ddr4_dqs_t,
  output [0:0]c1_ddr4_odt,
  output c1_ddr4_par,
  output c1_ddr4_reset_n,
  output c1_init_calib_complete,
  input  c0_init_calib_complete,
  input  c2_init_calib_complete,
  input  c3_init_calib_complete,
  output clk_out_125M,
  output clk_out_300M,
  output clk_out_400M,
  output clk_out_250M,
  output clk_out_PROG,
  input  MIG_1_RST,
  input sys_clk_gt,
  input sys_rst_n,
  input wire [1:0]cfg_current_speed,
  input wire cfg_err_cor_out,
  input wire cfg_err_fatal_out,
  input wire cfg_err_nonfatal_out,
  input wire [15:0]cfg_function_status,
  input wire [4:0]cfg_local_error_out,
  input wire [5:0]cfg_ltssm_state,
  input wire [1:0]cfg_max_payload,
  input wire [2:0]cfg_max_read_req,
  input wire [2:0]cfg_negotiated_width,
  input wire cfg_phy_link_down,
  input wire [1:0]cfg_phy_link_status,
  input wire cfg_pl_status_change,
  input wire [511:0]m_axis_cq_tdata,
  input wire [15:0]m_axis_cq_tkeep,
  input wire m_axis_cq_tlast,
  output wire m_axis_cq_tready,
  input wire [182:0]m_axis_cq_tuser,
  input wire m_axis_cq_tvalid,
  input wire [511:0]m_axis_rc_tdata,
  input wire [15:0]m_axis_rc_tkeep,
  input wire m_axis_rc_tlast,
  output wire m_axis_rc_tready,
  input wire [160:0]m_axis_rc_tuser,
  input wire m_axis_rc_tvalid,
  output wire [1:0]m_pcie_cq_np_req,
  output wire [7:0]pcie4_cfg_control_ds_bus_number,
  output wire [4:0]pcie4_cfg_control_ds_device_number,
  output wire [7:0]pcie4_cfg_control_ds_port_number,
  output wire [63:0]pcie4_cfg_control_dsn,
  output wire pcie4_cfg_control_err_cor_in,
  output wire pcie4_cfg_control_err_uncor_in,
  output wire [3:0]pcie4_cfg_control_flr_done,
  input wire [3:0]pcie4_cfg_control_flr_in_process,
  input wire pcie4_cfg_control_hot_reset_out,
  output wire pcie4_cfg_control_link_training_enable,
  input wire [251:0]pcie4_cfg_control_vf_flr_in_process,
  input wire [7:0]pcie4_cfg_fc_nph,
  output wire [2:0]pcie4_cfg_fc_sel,
  output wire [3:0]pcie4_cfg_interrupt_intx_vector,
  output wire [3:0]pcie4_cfg_interrupt_pending,
  input wire pcie4_cfg_interrupt_sent,
  input wire pcie4_cfg_mesg_rcvd_recd,
  input wire [7:0]pcie4_cfg_mesg_rcvd_recd_data,
  input wire [4:0]pcie4_cfg_mesg_rcvd_recd_type,
  output wire pcie4_cfg_mesg_tx_transmit,
  output wire [31:0]pcie4_cfg_mesg_tx_transmit_data,
  input wire pcie4_cfg_mesg_tx_transmit_done,
  output wire [2:0]pcie4_cfg_mesg_tx_transmit_type,
  output wire [9:0]pcie4_cfg_mgmt_addr,
  output wire [3:0]pcie4_cfg_mgmt_byte_en,
  output wire pcie4_cfg_mgmt_debug_access,
  output wire [7:0]pcie4_cfg_mgmt_function_number,
  input wire [31:0]pcie4_cfg_mgmt_read_data,
  output wire pcie4_cfg_mgmt_read_en,
  input wire pcie4_cfg_mgmt_read_write_done,
  output wire [31:0]pcie4_cfg_mgmt_write_data,
  output wire pcie4_cfg_mgmt_write_en,
  output wire [2:0]pcie4_cfg_msi_attr,
  input wire [31:0]pcie4_cfg_msi_data,
  input wire [3:0]pcie4_cfg_msi_enable,
  input wire pcie4_cfg_msi_fail,
  output wire [7:0]pcie4_cfg_msi_function_number,
  output wire [31:0]pcie4_cfg_msi_int_vector,
  input wire pcie4_cfg_msi_mask_update,
  output wire [31:0]pcie4_cfg_msi_pending_status,
  output wire pcie4_cfg_msi_pending_status_data_enable,
  output wire [3:0]pcie4_cfg_msi_pending_status_function_num,
  input wire pcie4_cfg_msi_sent,
  output wire pcie4_cfg_msi_tph_present,
  output wire [8:0]pcie4_cfg_msi_tph_st_tag,
  output wire [1:0]pcie4_cfg_msi_tph_type,
  input wire [5:0]pcie_cq_np_req_count,
  input wire [5:0]pcie_rq_seq_num0,
  input wire [5:0]pcie_rq_seq_num1,
  input wire pcie_rq_seq_num_vld0,
  input wire pcie_rq_seq_num_vld1,
  input wire phy_rdy_out,
  output wire [511:0]s_axis_cc_tdata,
  output wire [15:0]s_axis_cc_tkeep,
  output wire s_axis_cc_tlast,
  input wire s_axis_cc_tready,
  output wire [80:0]s_axis_cc_tuser,
  output wire s_axis_cc_tvalid,
  output wire [511:0]s_axis_rq_tdata,
  output wire [15:0]s_axis_rq_tkeep,
  output wire s_axis_rq_tlast,
  input wire [3:0]s_axis_rq_tready,
  output wire [136:0]s_axis_rq_tuser,
  output wire s_axis_rq_tvalid,
  input wire iiC_scl_i,
  output wire iiC_scl_o,
  output wire iiC_scl_t,
  input wire iiC_sda_i,
  output wire iiC_sda_o,
  output wire iiC_sda_t,
  input wire user_clk,
  input  wire user_lnk_up,
  input wire user_reset);

  wire [3:0]INIT_CAL_DONE;

  wire [31:0] EFUSE_IN_tri_i;
  reg [31:0] SHELL_VERSION_NUMBER = `SHELL_VERSION_NUMBER; // defined in shell_parameters.vh 

  wire [31:0]M_AXI_B_araddr;
  wire [2:0]M_AXI_B_arprot;
  wire M_AXI_B_arready;
  wire M_AXI_B_arvalid;
  wire [31:0]M_AXI_B_awaddr;
  wire [2:0]M_AXI_B_awprot;
  wire M_AXI_B_awready;
  wire M_AXI_B_awvalid;
  wire M_AXI_B_bready;
  wire [1:0]M_AXI_B_bresp;
  wire M_AXI_B_bvalid;
  wire [31:0]M_AXI_B_rdata;
  wire M_AXI_B_rready;
  wire [1:0]M_AXI_B_rresp;
  wire M_AXI_B_rvalid;
  wire [31:0]M_AXI_B_wdata;
  wire M_AXI_B_wready;
  wire [3:0]M_AXI_B_wstrb;
  wire M_AXI_B_wvalid;

  wire clk_250M;

  wire axi_aresetn;

  assign EFUSE_IN_tri_i =  32'h12345566;

  assign INIT_CAL_DONE = {c0_init_calib_complete, c1_init_calib_complete, c2_init_calib_complete, c3_init_calib_complete};

  assign clk_out_250M = clk_250M;


  PL_X PL_X_i
       (.BMC_GPIO(BMC_GPIO),
        .BMC_UART_rxd(BMC_UART_rxd),
        .BMC_UART_txd(BMC_UART_txd),
        .C0_DDR_SREF_CTRL_IN(C0_DDR_SREF_CTRL_IN),
        .C0_DDR_SREF_CTRL_OUT(C0_DDR_SREF_CTRL_OUT),
        .C1_SYS_CLK(C1_SYS_CLK),
        .C2_DDR_SREF_CTRL_IN(C2_DDR_SREF_CTRL_IN),
        .C2_DDR_SREF_CTRL_OUT(C2_DDR_SREF_CTRL_OUT),
        .C3_DDR_SREF_CTRL_IN(C3_DDR_SREF_CTRL_IN),
        .C3_DDR_SREF_CTRL_OUT(C3_DDR_SREF_CTRL_OUT),
        .EFUSE_IN_tri_i(EFUSE_IN_tri_i),
        .INIT_CAL_DONE(INIT_CAL_DONE),
        .MIG_1_RST(MIG_1_RST),
        .M_AXI_LITE_TO_HLS_PR_NORTH_araddr(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_araddr),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arprot(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arprot),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awaddr(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awaddr),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awprot(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awprot),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bresp(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bresp),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rdata(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rdata),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rresp(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rresp),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wdata(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wdata),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wstrb(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wstrb),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wvalid),
        .S00_AXI_0_araddr(M_AXI_B_araddr),
        .S00_AXI_0_arprot(M_AXI_B_arprot),
        .S00_AXI_0_arready(M_AXI_B_arready),
        .S00_AXI_0_arvalid(M_AXI_B_arvalid),
        .S00_AXI_0_awaddr(M_AXI_B_awaddr),
        .S00_AXI_0_awprot(M_AXI_B_awprot),
        .S00_AXI_0_awready(M_AXI_B_awready),
        .S00_AXI_0_awvalid(M_AXI_B_awvalid),
        .S00_AXI_0_bready(M_AXI_B_bready),
        .S00_AXI_0_bresp(M_AXI_B_bresp),
        .S00_AXI_0_bvalid(M_AXI_B_bvalid),
        .S00_AXI_0_rdata(M_AXI_B_rdata),
        .S00_AXI_0_rready(M_AXI_B_rready),
        .S00_AXI_0_rresp(M_AXI_B_rresp),
        .S00_AXI_0_rvalid(M_AXI_B_rvalid),
        .S00_AXI_0_wdata(M_AXI_B_wdata),
        .S00_AXI_0_wready(M_AXI_B_wready),
        .S00_AXI_0_wstrb(M_AXI_B_wstrb),
        .S00_AXI_0_wvalid(M_AXI_B_wvalid),
        .SHELL_VERSION_IN_tri_i(SHELL_VERSION_NUMBER),
        .S_AXI_MM_0_araddr(S_AXI_MM_MIG.AXI_araddr),
        .S_AXI_MM_0_arburst(S_AXI_MM_MIG.AXI_arburst),
        .S_AXI_MM_0_arcache(S_AXI_MM_MIG.AXI_arcache),
        .S_AXI_MM_0_arid(S_AXI_MM_MIG.AXI_arid),
        .S_AXI_MM_0_arlen(S_AXI_MM_MIG.AXI_arlen),
        .S_AXI_MM_0_arlock(S_AXI_MM_MIG.AXI_arlock),
        .S_AXI_MM_0_arprot(S_AXI_MM_MIG.AXI_arprot),
        .S_AXI_MM_0_arqos(S_AXI_MM_MIG.AXI_arqos),
        .S_AXI_MM_0_arready(S_AXI_MM_MIG.AXI_arready),
        .S_AXI_MM_0_arregion(S_AXI_MM_MIG.AXI_arregion),
        .S_AXI_MM_0_arsize(S_AXI_MM_MIG.AXI_arsize),
        .S_AXI_MM_0_arvalid(S_AXI_MM_MIG.AXI_arvalid),
        .S_AXI_MM_0_awaddr(S_AXI_MM_MIG.AXI_awaddr),
        .S_AXI_MM_0_awburst(S_AXI_MM_MIG.AXI_awburst),
        .S_AXI_MM_0_awcache(S_AXI_MM_MIG.AXI_awcache),
        .S_AXI_MM_0_awid(S_AXI_MM_MIG.AXI_awid),
        .S_AXI_MM_0_awlen(S_AXI_MM_MIG.AXI_awlen),
        .S_AXI_MM_0_awlock(S_AXI_MM_MIG.AXI_awlock),
        .S_AXI_MM_0_awprot(S_AXI_MM_MIG.AXI_awprot),
        .S_AXI_MM_0_awqos(S_AXI_MM_MIG.AXI_awqos),
        .S_AXI_MM_0_awready(S_AXI_MM_MIG.AXI_awready),
        .S_AXI_MM_0_awregion(S_AXI_MM_MIG.AXI_awregion),
        .S_AXI_MM_0_awsize(S_AXI_MM_MIG.AXI_awsize),
        .S_AXI_MM_0_awvalid(S_AXI_MM_MIG.AXI_awvalid),
        .S_AXI_MM_0_bid(S_AXI_MM_MIG.AXI_bid),
        .S_AXI_MM_0_bready(S_AXI_MM_MIG.AXI_bready),
        .S_AXI_MM_0_bresp(S_AXI_MM_MIG.AXI_bresp),
        .S_AXI_MM_0_bvalid(S_AXI_MM_MIG.AXI_bvalid),
        .S_AXI_MM_0_rdata(S_AXI_MM_MIG.AXI_rdata),
        .S_AXI_MM_0_rid(S_AXI_MM_MIG.AXI_rid),
        .S_AXI_MM_0_rlast(S_AXI_MM_MIG.AXI_rlast),
        .S_AXI_MM_0_rready(S_AXI_MM_MIG.AXI_rready),
        .S_AXI_MM_0_rresp(S_AXI_MM_MIG.AXI_rresp),
        .S_AXI_MM_0_rvalid(S_AXI_MM_MIG.AXI_rvalid),
        .S_AXI_MM_0_wdata(S_AXI_MM_MIG.AXI_wdata),
        .S_AXI_MM_0_wlast(S_AXI_MM_MIG.AXI_wlast),
        .S_AXI_MM_0_wready(S_AXI_MM_MIG.AXI_wready),
        .S_AXI_MM_0_wstrb(S_AXI_MM_MIG.AXI_wstrb),
        .S_AXI_MM_0_wvalid(S_AXI_MM_MIG.AXI_wvalid),
        .axi_reset_n_250M_out(axi_reset_n_out),
        .c1_ddr4_act_n(c1_ddr4_act_n),
        .c1_ddr4_adr(c1_ddr4_adr),
        .c1_ddr4_ba(c1_ddr4_ba),
        .c1_ddr4_bg(c1_ddr4_bg),
        .c1_ddr4_ck_c(c1_ddr4_ck_c),
        .c1_ddr4_ck_t(c1_ddr4_ck_t),
        .c1_ddr4_cke(c1_ddr4_cke),
        .c1_ddr4_cs_n(c1_ddr4_cs_n),
        .c1_ddr4_dq(c1_ddr4_dq),
        .c1_ddr4_dqs_c(c1_ddr4_dqs_c),
        .c1_ddr4_dqs_t(c1_ddr4_dqs_t),
        .c1_ddr4_odt(c1_ddr4_odt),
        .c1_ddr4_par(c1_ddr4_par),
        .c1_ddr4_reset_n(c1_ddr4_reset_n),
        .c1_init_calib_complete(c1_init_calib_complete),
        .clk_250M(clk_250M),
        .clk_out_125M(clk_out_125M),
        .clk_out_300M(clk_out_300M),
        .clk_out_400M(clk_out_400M),
        .clk_out_PROG(clk_out_PROG),
        .deviceDNA_PA_tri_i(32'h12345678),
        .deviceDNA_PB_tri_i(32'hABCDEF00),
        .deviceDNA_PC_tri_i(32'hFEEDBEEF),
        .deviceDNA_PD_tri_i(32'haa556699),
        .iiC_scl_i(iiC_scl_i),
        .iiC_scl_o(iiC_scl_o),
        .iiC_scl_t(iiC_scl_t),
        .iiC_sda_i(iiC_sda_i),
        .iiC_sda_o(iiC_sda_o),
        .iiC_sda_t(iiC_sda_t),
        .s_axi_aresetn(axi_aresetn),
        .user_lnk_up_sd(user_lnk_up));


  X_PCIe_Bridge_ICAP_complex PCIe_Bridge_ICAP_complex_i (
        .M_AXI_B_araddr(M_AXI_B_araddr),
        .M_AXI_B_arprot(M_AXI_B_arprot),
        .M_AXI_B_arready(M_AXI_B_arready),
        .M_AXI_B_aruser(),
        .M_AXI_B_arvalid(M_AXI_B_arvalid),
        .M_AXI_B_awaddr(M_AXI_B_awaddr),
        .M_AXI_B_awprot(M_AXI_B_awprot),
        .M_AXI_B_awready(M_AXI_B_awready),
        .M_AXI_B_awuser(),
        .M_AXI_B_awvalid(M_AXI_B_awvalid),
        .M_AXI_B_bready(M_AXI_B_bready),
        .M_AXI_B_bresp(M_AXI_B_bresp),
        .M_AXI_B_bvalid(M_AXI_B_bvalid),
        .M_AXI_B_rdata(M_AXI_B_rdata),
        .M_AXI_B_rready(M_AXI_B_rready),
        .M_AXI_B_rresp(M_AXI_B_rresp),
        .M_AXI_B_rvalid(M_AXI_B_rvalid),
        .M_AXI_B_wdata(M_AXI_B_wdata),
        .M_AXI_B_wready(M_AXI_B_wready),
        .M_AXI_B_wstrb(M_AXI_B_wstrb),
        .M_AXI_B_wvalid(M_AXI_B_wvalid),
        .S_AXI_MM_PCIM_araddr(S_AXI_MM_PCIM.AXI_araddr),
        .S_AXI_MM_PCIM_arburst(S_AXI_MM_PCIM.AXI_arburst),
        .S_AXI_MM_PCIM_arid(S_AXI_MM_PCIM.AXI_arid),
        .S_AXI_MM_PCIM_arlen(S_AXI_MM_PCIM.AXI_arlen),
        .S_AXI_MM_PCIM_arready(S_AXI_MM_PCIM.AXI_arready),
        .S_AXI_MM_PCIM_arregion(S_AXI_MM_PCIM.AXI_arregion),
        .S_AXI_MM_PCIM_arsize(S_AXI_MM_PCIM.AXI_arsize),
        .S_AXI_MM_PCIM_arvalid(S_AXI_MM_PCIM.AXI_arvalid),
        .S_AXI_MM_PCIM_awaddr(S_AXI_MM_PCIM.AXI_awaddr),
        .S_AXI_MM_PCIM_awburst(S_AXI_MM_PCIM.AXI_awburst),
        .S_AXI_MM_PCIM_awid(S_AXI_MM_PCIM.AXI_awid),
        .S_AXI_MM_PCIM_awlen(S_AXI_MM_PCIM.AXI_awlen),
        .S_AXI_MM_PCIM_awready(S_AXI_MM_PCIM.AXI_awready),
        .S_AXI_MM_PCIM_awregion(S_AXI_MM_PCIM.AXI_awregion),
        .S_AXI_MM_PCIM_awsize(S_AXI_MM_PCIM.AXI_awsize),
        .S_AXI_MM_PCIM_awvalid(S_AXI_MM_PCIM.AXI_awvalid),
        .S_AXI_MM_PCIM_bid(S_AXI_MM_PCIM.AXI_bid),
        .S_AXI_MM_PCIM_bready(S_AXI_MM_PCIM.AXI_bready),
        .S_AXI_MM_PCIM_bresp(S_AXI_MM_PCIM.AXI_bresp),
        .S_AXI_MM_PCIM_bvalid(S_AXI_MM_PCIM.AXI_bvalid),
        .S_AXI_MM_PCIM_rdata(S_AXI_MM_PCIM.AXI_rdata),
        .S_AXI_MM_PCIM_rid(S_AXI_MM_PCIM.AXI_rid),
        .S_AXI_MM_PCIM_rlast(S_AXI_MM_PCIM.AXI_rlast),
        .S_AXI_MM_PCIM_rready(S_AXI_MM_PCIM.AXI_rready),
        .S_AXI_MM_PCIM_rresp(S_AXI_MM_PCIM.AXI_rresp),
        .S_AXI_MM_PCIM_ruser(),
        .S_AXI_MM_PCIM_rvalid(S_AXI_MM_PCIM.AXI_rvalid),
        .S_AXI_MM_PCIM_wdata(S_AXI_MM_PCIM.AXI_wdata),
        .S_AXI_MM_PCIM_wlast(S_AXI_MM_PCIM.AXI_wlast),
        .S_AXI_MM_PCIM_wready(S_AXI_MM_PCIM.AXI_wready),
        .S_AXI_MM_PCIM_wstrb(S_AXI_MM_PCIM.AXI_wstrb),
        .S_AXI_MM_PCIM_wuser(64'd0),
        .S_AXI_MM_PCIM_wvalid(S_AXI_MM_PCIM.AXI_wvalid),
        .axi_aresetn(axi_aresetn),
        .clk_out_250M(clk_250M),
        .sys_rst_n(sys_rst_n),
  .cfg_current_speed(cfg_current_speed),
  .cfg_err_cor_out(cfg_err_cor_out),
  .cfg_err_fatal_out(cfg_err_fatal_out),
  .cfg_err_nonfatal_out(cfg_err_nonfatal_out),
  .cfg_function_status(cfg_function_status),
  .cfg_local_error_out(cfg_local_error_out),
  .cfg_ltssm_state(cfg_ltssm_state),
  .cfg_max_payload(cfg_max_payload),
  .cfg_max_read_req(cfg_max_read_req),
  .cfg_negotiated_width(cfg_negotiated_width),
  .cfg_phy_link_down(cfg_phy_link_down),
  .cfg_phy_link_status(cfg_phy_link_status),
  .cfg_pl_status_change(cfg_pl_status_change),
  .m_axis_cq_tdata(m_axis_cq_tdata),
  .m_axis_cq_tkeep(m_axis_cq_tkeep),
  .m_axis_cq_tlast(m_axis_cq_tlast),
  .m_axis_cq_tready(m_axis_cq_tready),
  .m_axis_cq_tuser(m_axis_cq_tuser),
  .m_axis_cq_tvalid(m_axis_cq_tvalid),
  .m_axis_rc_tdata(m_axis_rc_tdata),
  .m_axis_rc_tkeep(m_axis_rc_tkeep),
  .m_axis_rc_tlast(m_axis_rc_tlast),
  .m_axis_rc_tready(m_axis_rc_tready),
  .m_axis_rc_tuser(m_axis_rc_tuser),
  .m_axis_rc_tvalid(m_axis_rc_tvalid),
  .m_pcie_cq_np_req(m_pcie_cq_np_req),
  .pcie4_cfg_control_ds_bus_number(pcie4_cfg_control_ds_bus_number),
  .pcie4_cfg_control_ds_device_number(pcie4_cfg_control_ds_device_number),
  .pcie4_cfg_control_ds_port_number(pcie4_cfg_control_ds_port_number),
  .pcie4_cfg_control_dsn(pcie4_cfg_control_dsn),
  .pcie4_cfg_control_err_cor_in(pcie4_cfg_control_err_cor_in),
  .pcie4_cfg_control_err_uncor_in(pcie4_cfg_control_err_uncor_in),
  .pcie4_cfg_control_flr_done(pcie4_cfg_control_flr_done),
  .pcie4_cfg_control_flr_in_process(pcie4_cfg_control_flr_in_process),
  .pcie4_cfg_control_hot_reset_out(pcie4_cfg_control_hot_reset_out),
  .pcie4_cfg_control_link_training_enable(pcie4_cfg_control_link_training_enable),
  .pcie4_cfg_control_vf_flr_in_process(pcie4_cfg_control_vf_flr_in_process),
  .pcie4_cfg_fc_nph(pcie4_cfg_fc_nph),
  .pcie4_cfg_fc_sel(pcie4_cfg_fc_sel),
  .pcie4_cfg_interrupt_intx_vector(pcie4_cfg_interrupt_intx_vector),
  .pcie4_cfg_interrupt_pending(pcie4_cfg_interrupt_pending),
  .pcie4_cfg_interrupt_sent(pcie4_cfg_interrupt_sent),
  .pcie4_cfg_mesg_rcvd_recd(pcie4_cfg_mesg_rcvd_recd),
  .pcie4_cfg_mesg_rcvd_recd_data(pcie4_cfg_mesg_rcvd_recd_data),
  .pcie4_cfg_mesg_rcvd_recd_type(pcie4_cfg_mesg_rcvd_recd_type),
  .pcie4_cfg_mesg_tx_transmit(pcie4_cfg_mesg_tx_transmit),
  .pcie4_cfg_mesg_tx_transmit_data(pcie4_cfg_mesg_tx_transmit_data),
  .pcie4_cfg_mesg_tx_transmit_done(pcie4_cfg_mesg_tx_transmit_done),
  .pcie4_cfg_mesg_tx_transmit_type(pcie4_cfg_mesg_tx_transmit_type),
  .pcie4_cfg_mgmt_addr(pcie4_cfg_mgmt_addr),
  .pcie4_cfg_mgmt_byte_en(pcie4_cfg_mgmt_byte_en),
  .pcie4_cfg_mgmt_debug_access(pcie4_cfg_mgmt_debug_access),
  .pcie4_cfg_mgmt_function_number(pcie4_cfg_mgmt_function_number),
  .pcie4_cfg_mgmt_read_data(pcie4_cfg_mgmt_read_data),
  .pcie4_cfg_mgmt_read_en(pcie4_cfg_mgmt_read_en),
  .pcie4_cfg_mgmt_read_write_done(pcie4_cfg_mgmt_read_write_done),
  .pcie4_cfg_mgmt_write_data(pcie4_cfg_mgmt_write_data),
  .pcie4_cfg_mgmt_write_en(pcie4_cfg_mgmt_write_en),
  .pcie4_cfg_msi_attr(pcie4_cfg_msi_attr),
  .pcie4_cfg_msi_data(pcie4_cfg_msi_data),
  .pcie4_cfg_msi_enable(pcie4_cfg_msi_enable),
  .pcie4_cfg_msi_fail(pcie4_cfg_msi_fail),
  .pcie4_cfg_msi_function_number(pcie4_cfg_msi_function_number),
  .pcie4_cfg_msi_int_vector(pcie4_cfg_msi_int_vector),
  .pcie4_cfg_msi_mask_update(pcie4_cfg_msi_mask_update),
  .pcie4_cfg_msi_pending_status(pcie4_cfg_msi_pending_status),
  .pcie4_cfg_msi_pending_status_data_enable(pcie4_cfg_msi_pending_status_data_enable),
  .pcie4_cfg_msi_pending_status_function_num(pcie4_cfg_msi_pending_status_function_num),
  .pcie4_cfg_msi_sent(pcie4_cfg_msi_sent),
  .pcie4_cfg_msi_tph_present(pcie4_cfg_msi_tph_present),
  .pcie4_cfg_msi_tph_st_tag(pcie4_cfg_msi_tph_st_tag),
  .pcie4_cfg_msi_tph_type(pcie4_cfg_msi_tph_type),
  .pcie_cq_np_req_count(pcie_cq_np_req_count),
  .pcie_rq_seq_num0(pcie_rq_seq_num0),
  .pcie_rq_seq_num1(pcie_rq_seq_num1),
  .pcie_rq_seq_num_vld0(pcie_rq_seq_num_vld0),
  .pcie_rq_seq_num_vld1(pcie_rq_seq_num_vld1),
  .phy_rdy_out(phy_rdy_out),
  .s_axis_cc_tdata(s_axis_cc_tdata),
  .s_axis_cc_tkeep(s_axis_cc_tkeep),
  .s_axis_cc_tlast(s_axis_cc_tlast),
  .s_axis_cc_tready(s_axis_cc_tready),
  .s_axis_cc_tuser(s_axis_cc_tuser),
  .s_axis_cc_tvalid(s_axis_cc_tvalid),
  .s_axis_rq_tdata(s_axis_rq_tdata),
  .s_axis_rq_tkeep(s_axis_rq_tkeep),
  .s_axis_rq_tlast(s_axis_rq_tlast),
  .s_axis_rq_tready(s_axis_rq_tready),
  .s_axis_rq_tuser(s_axis_rq_tuser),
  .s_axis_rq_tvalid(s_axis_rq_tvalid),
  .user_clk(user_clk),
  .user_lnk_up(user_lnk_up),
  .user_reset(user_reset));


endmodule
